
//=========================== All Files ===============================
//----> Impoting the package
`include "uvm_pkg.sv"
import uvm_pkg::*;

//----> Including the files
`include "fa_common.sv"
`include "full_adder.v"
`include "fa_inf.sv"
`include "fa_tx.sv"
`include "fa_seq_lib.sv"
`include "fa_sqr.sv"
`include "fa_driver.sv"
`include "fa_monitor.sv"
`include "fa_coverage.sv"
`include "fa_agent.sv"
`include "fa_scoreboard.sv"
`include "fa_env.sv"
`include "fa_test_lib.sv"
`include "top.sv"

//======================================================================
// This file includes all the files required for the full adder testbench

