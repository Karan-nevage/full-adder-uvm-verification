// ======================== Full Adder Sequencer ==================================

class fa_sqr extends uvm_sequencer#(fa_tx);
    `uvm_component_utils(fa_sqr)
    `NEW_COMP
endclass

//===============================================================================
// This file contains the sequencer for the full adder component