// ========================= Full Adder Interface ==============================  

interface fa_intf();
    logic a;
    logic b;
    logic cin;
    logic sum;
    logic cout;
endinterface

//===============================================================================
// This file contains the interface for the full adder component